2
2 2 2 2 2 r h 46 B 0 B
2 2 2 2 2 r h 8 B 50 H
20 20 20 20 20 r 53 57 58 65 h 27 T 52 T 20 T
3 3 3 3 3 r h 44 T 32 B
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
5
