3
0 0 0 0 0 r 18 22 h 37 B 25 B 13 B
1 3 1 0 2 r 61 57 h 44 T 32 H 20 B
20 17 15 8 25 r 23 32 h 39 T 27 T 15 T
90 90 90 90 90 r 33 41 h 46 T 34 H 22 B
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
9
